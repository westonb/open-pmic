magic
tech sky130A
magscale 1 2
timestamp 1618785568
<< error_p >>
rect -410 660 -394 676
rect 394 660 410 676
rect -426 644 -410 660
rect 410 644 426 660
rect -426 620 -410 636
rect 410 620 426 636
rect -410 604 -394 620
rect 394 604 410 620
rect -660 410 -644 426
rect -636 410 -620 426
rect 620 410 636 426
rect 644 410 660 426
rect -676 394 -660 410
rect -620 394 -604 410
rect 604 394 620 410
rect 660 394 676 410
rect -676 -410 -660 -394
rect -620 -410 -604 -394
rect 604 -410 620 -394
rect 660 -410 676 -394
rect -660 -426 -644 -410
rect -636 -426 -620 -410
rect 620 -426 636 -410
rect 644 -426 660 -410
rect -410 -620 -394 -604
rect 394 -620 410 -604
rect -426 -636 -410 -620
rect 410 -636 426 -620
rect -426 -660 -410 -644
rect 410 -660 426 -644
rect -410 -676 -394 -660
rect 394 -676 410 -660
<< mvnmos >>
rect -460 500 460 600
rect -600 -460 -500 460
rect 500 -460 600 460
rect -460 -600 460 -500
<< mvndiff >>
rect -700 680 -400 700
rect 400 680 700 700
rect -700 660 700 680
rect -700 640 -410 660
rect -700 460 -640 640
rect -460 620 -410 640
rect 410 640 700 660
rect 410 620 460 640
rect -460 600 460 620
rect -460 480 460 500
rect -460 460 -410 480
rect -700 410 -600 460
rect -700 400 -660 410
rect -680 -400 -660 400
rect -700 -410 -660 -400
rect -620 -410 -600 410
rect -700 -460 -600 -410
rect -500 440 -410 460
rect 410 460 460 480
rect 640 460 700 640
rect 410 440 500 460
rect -500 420 500 440
rect -500 410 -400 420
rect -500 -410 -480 410
rect -440 400 -400 410
rect 400 410 500 420
rect 400 400 440 410
rect -440 -400 -420 400
rect 420 -400 440 400
rect -440 -410 -400 -400
rect -500 -420 -400 -410
rect 400 -410 440 -400
rect 480 -410 500 410
rect 400 -420 500 -410
rect -500 -440 500 -420
rect -500 -460 -410 -440
rect -700 -640 -640 -460
rect -460 -480 -410 -460
rect 410 -460 500 -440
rect 600 410 700 460
rect 600 -410 620 410
rect 660 400 700 410
rect 660 -400 680 400
rect 660 -410 700 -400
rect 600 -460 700 -410
rect 410 -480 460 -460
rect -460 -500 460 -480
rect -460 -620 460 -600
rect -460 -640 -410 -620
rect -700 -660 -410 -640
rect 410 -640 460 -620
rect 640 -640 700 -460
rect 410 -660 700 -640
rect -700 -680 700 -660
rect -700 -700 -410 -680
rect 400 -700 700 -680
<< mvndiffc >>
rect -410 620 410 660
rect -660 -410 -620 410
rect -410 440 410 480
rect -480 -410 -440 410
rect 440 -410 480 410
rect -410 -480 410 -440
rect 620 -410 660 410
rect -410 -660 410 -620
<< poly >>
rect -600 580 -460 600
rect -600 520 -580 580
rect -520 520 -460 580
rect -600 500 -460 520
rect 460 580 600 600
rect 460 520 520 580
rect 580 520 600 580
rect 460 500 600 520
rect -600 460 -500 500
rect 500 460 600 500
rect -600 -500 -500 -460
rect 500 -500 600 -460
rect -600 -520 -460 -500
rect -600 -580 -580 -520
rect -520 -580 -460 -520
rect -600 -600 -460 -580
rect 460 -520 600 -500
rect 460 -580 520 -520
rect 580 -580 600 -520
rect 460 -600 600 -580
<< polycont >>
rect -580 520 -520 580
rect 520 520 580 580
rect -580 -580 -520 -520
rect 520 -580 580 -520
<< locali >>
rect -600 580 -500 600
rect -600 520 -580 580
rect -520 520 -500 580
rect -600 500 -500 520
rect 500 580 600 600
rect 500 520 520 580
rect 580 520 600 580
rect 500 500 600 520
rect -460 460 -410 480
rect -480 440 -410 460
rect 410 460 460 480
rect 410 440 480 460
rect -480 430 -400 440
rect 400 430 480 440
rect -480 420 480 430
rect -480 410 -420 420
rect -440 400 -420 410
rect -430 -400 -420 400
rect -440 -410 -420 -400
rect -480 -420 -420 -410
rect 420 410 480 420
rect 420 400 440 410
rect 420 -400 430 400
rect 420 -410 440 -400
rect 420 -420 480 -410
rect -480 -430 480 -420
rect -480 -440 -400 -430
rect 400 -440 480 -430
rect -480 -460 -410 -440
rect -460 -480 -410 -460
rect 410 -460 480 -440
rect 410 -480 460 -460
rect -600 -520 -500 -500
rect -600 -580 -580 -520
rect -520 -580 -500 -520
rect -600 -600 -500 -580
rect 500 -520 600 -500
rect 500 -580 520 -520
rect 580 -580 600 -520
rect 500 -600 600 -580
<< viali >>
rect -580 520 -520 580
rect 520 520 580 580
rect -400 440 400 470
rect -400 430 400 440
rect -470 -400 -440 400
rect -440 -400 -430 400
rect 430 -400 440 400
rect 440 -400 470 400
rect -400 -440 400 -430
rect -400 -470 400 -440
rect -580 -580 -520 -520
rect 520 -580 580 -520
<< metal1 >>
rect -600 580 -500 600
rect -600 520 -580 580
rect -520 520 -500 580
rect -600 500 -500 520
rect 500 580 600 600
rect 500 520 520 580
rect 580 520 600 580
rect 500 500 600 520
rect -440 470 440 480
rect -440 440 -400 470
rect -480 430 -400 440
rect 400 440 440 470
rect 400 430 480 440
rect -480 400 480 430
rect -480 -400 -470 400
rect -430 280 430 400
rect -430 200 -280 280
rect -200 200 -160 280
rect -80 200 -40 280
rect 40 200 80 280
rect 160 200 430 280
rect -430 160 430 200
rect -430 80 -280 160
rect -200 80 -160 160
rect -80 80 -40 160
rect 40 80 80 160
rect 160 80 200 160
rect 280 80 430 160
rect -430 40 430 80
rect -430 -40 -280 40
rect -200 -40 -160 40
rect -80 -40 -40 40
rect 40 -40 80 40
rect 160 -40 200 40
rect 280 -40 430 40
rect -430 -80 430 -40
rect -430 -160 -280 -80
rect -200 -160 -160 -80
rect -80 -160 -40 -80
rect 40 -160 80 -80
rect 160 -160 200 -80
rect 280 -160 430 -80
rect -430 -200 430 -160
rect -430 -280 -160 -200
rect -80 -280 -40 -200
rect 40 -280 80 -200
rect 160 -280 200 -200
rect 280 -280 430 -200
rect -430 -400 430 -280
rect 470 -400 480 400
rect -480 -430 480 -400
rect -480 -440 -400 -430
rect -440 -470 -400 -440
rect 400 -440 480 -430
rect 400 -470 440 -440
rect -440 -480 440 -470
rect -600 -520 -500 -500
rect -600 -580 -580 -520
rect -520 -580 -500 -520
rect -600 -600 -500 -580
rect 500 -520 600 -500
rect 500 -580 520 -520
rect 580 -580 600 -520
rect 500 -600 600 -580
<< via1 >>
rect -580 520 -520 580
rect 520 520 580 580
rect -280 200 -200 280
rect -160 200 -80 280
rect -40 200 40 280
rect 80 200 160 280
rect -280 80 -200 160
rect -160 80 -80 160
rect -40 80 40 160
rect 80 80 160 160
rect 200 80 280 160
rect -280 -40 -200 40
rect -160 -40 -80 40
rect -40 -40 40 40
rect 80 -40 160 40
rect 200 -40 280 40
rect -280 -160 -200 -80
rect -160 -160 -80 -80
rect -40 -160 40 -80
rect 80 -160 160 -80
rect 200 -160 280 -80
rect -160 -280 -80 -200
rect -40 -280 40 -200
rect 80 -280 160 -200
rect 200 -280 280 -200
rect -580 -580 -520 -520
rect 520 -580 580 -520
<< metal2 >>
rect -600 580 600 600
rect -600 520 -580 580
rect -520 520 520 580
rect 580 520 600 580
rect -600 500 600 520
rect -600 -500 -500 500
rect -400 280 80 400
tri 80 280 200 400 sw
rect -400 200 -280 280
rect -200 200 -160 280
rect -80 200 -40 280
rect 40 200 80 280
rect 160 200 200 280
rect -400 160 200 200
tri 200 160 320 280 sw
rect -400 80 -280 160
rect -200 80 -160 160
rect -80 80 -40 160
rect 40 80 80 160
rect 160 80 200 160
rect 280 80 320 160
tri 320 80 400 160 sw
rect -400 40 400 80
rect -400 -40 -280 40
rect -200 -40 -160 40
rect -80 -40 -40 40
rect 40 -40 80 40
rect 160 -40 200 40
rect 280 -40 400 40
rect -400 -80 400 -40
tri -400 -200 -280 -80 ne
rect -200 -160 -160 -80
rect -80 -160 -40 -80
rect 40 -160 80 -80
rect 160 -160 200 -80
rect 280 -160 400 -80
rect -280 -200 400 -160
tri -280 -280 -200 -200 ne
rect -200 -280 -160 -200
rect -80 -280 -40 -200
rect 40 -280 80 -200
rect 160 -280 200 -200
rect 280 -280 400 -200
tri -200 -400 -80 -280 ne
rect -80 -400 400 -280
rect 500 -500 600 500
rect -600 -520 600 -500
rect -600 -580 -580 -520
rect -520 -580 520 -520
rect 580 -580 600 -520
rect -600 -600 600 -580
<< via2 >>
rect -280 200 -200 280
rect -160 200 -80 280
rect -40 200 40 280
rect 80 200 160 280
rect -280 80 -200 160
rect -160 80 -80 160
rect -40 80 40 160
rect 80 80 160 160
rect 200 80 280 160
rect -280 -40 -200 40
rect -160 -40 -80 40
rect -40 -40 40 40
rect 80 -40 160 40
rect 200 -40 280 40
rect -280 -160 -200 -80
rect -160 -160 -80 -80
rect -40 -160 40 -80
rect 80 -160 160 -80
rect 200 -160 280 -80
rect -160 -280 -80 -200
rect -40 -280 40 -200
rect 80 -280 160 -200
rect 200 -280 280 -200
<< metal3 >>
tri -1031 550 -550 1031 se
tri -1031 69 -550 550 ne
tri -550 280 201 1031 sw
rect -550 200 -280 280
rect -200 200 -160 280
rect -80 200 -40 280
rect 40 200 80 280
rect 160 200 201 280
rect -550 160 201 200
tri 201 160 321 280 sw
rect -550 80 -280 160
rect -200 80 -160 160
rect -80 80 -40 160
rect 40 80 80 160
rect 160 80 200 160
rect 280 80 321 160
rect -550 69 321 80
tri -550 -200 -281 69 ne
rect -281 40 321 69
rect -281 -40 -280 40
rect -200 -40 -160 40
rect -80 -40 -40 40
rect 40 -40 80 40
rect 160 -40 200 40
rect 280 -40 321 40
rect -281 -80 321 -40
tri 321 -80 561 160 sw
rect -281 -160 -280 -80
rect -200 -160 -160 -80
rect -80 -160 -40 -80
rect 40 -160 80 -80
rect 160 -160 200 -80
rect 280 -160 561 -80
rect -281 -200 561 -160
tri -281 -280 -201 -200 ne
rect -201 -280 -160 -200
rect -80 -280 -40 -200
rect 40 -280 80 -200
rect 160 -280 200 -200
rect 280 -280 561 -200
tri -201 -1031 550 -280 ne
rect 550 -550 561 -280
tri 561 -550 1031 -80 sw
tri 550 -1031 1031 -550 nw
<< via3 >>
rect -280 200 -200 280
rect -160 200 -80 280
rect -40 200 40 280
rect 80 200 160 280
rect -280 80 -200 160
rect -160 80 -80 160
rect -40 80 40 160
rect 80 80 160 160
rect 200 80 280 160
rect -280 -40 -200 40
rect -160 -40 -80 40
rect -40 -40 40 40
rect 80 -40 160 40
rect 200 -40 280 40
rect -280 -160 -200 -80
rect -160 -160 -80 -80
rect -40 -160 40 -80
rect 80 -160 160 -80
rect 200 -160 280 -80
rect -160 -280 -80 -200
rect -40 -280 40 -200
rect 80 -280 160 -200
rect 200 -280 280 -200
<< metal4 >>
tri -1031 550 -550 1031 se
tri -1031 69 -550 550 ne
tri -550 420 61 1031 sw
rect -550 180 -420 420
rect -180 280 61 420
tri 61 280 201 420 sw
rect -180 200 -160 280
rect -80 200 -40 280
rect 40 200 80 280
rect 160 200 201 280
rect -180 180 201 200
rect -550 160 201 180
tri 201 160 321 280 sw
rect -550 80 -280 160
rect -200 80 -160 160
rect -80 120 -40 160
rect 40 120 80 160
rect 160 80 200 160
rect 280 80 321 160
rect -550 69 -120 80
tri -550 -200 -281 69 ne
rect -281 40 -120 69
rect 120 50 321 80
tri 321 50 431 160 sw
rect 120 40 431 50
rect -281 -40 -280 40
rect -200 -40 -160 40
rect 160 -40 200 40
rect 280 -40 431 40
rect -281 -80 -120 -40
rect 120 -80 431 -40
rect -281 -160 -280 -80
rect -200 -160 -160 -80
rect -80 -160 -40 -120
rect 40 -160 80 -120
rect 160 -160 200 -80
rect 280 -160 431 -80
rect -281 -180 431 -160
rect -281 -200 180 -180
tri -281 -280 -201 -200 ne
rect -201 -280 -160 -200
rect -80 -280 -40 -200
rect 40 -280 80 -200
rect 160 -280 180 -200
tri -201 -550 69 -280 ne
rect 69 -420 180 -280
rect 420 -420 431 -180
rect 69 -550 431 -420
tri 431 -550 1031 50 sw
tri 69 -1031 550 -550 ne
tri 550 -1031 1031 -550 nw
<< via4 >>
rect -420 280 -180 420
rect -420 200 -280 280
rect -280 200 -200 280
rect -200 200 -180 280
rect -420 180 -180 200
rect -120 80 -80 120
rect -80 80 -40 120
rect -40 80 40 120
rect 40 80 80 120
rect 80 80 120 120
rect -120 40 120 80
rect -120 -40 -80 40
rect -80 -40 -40 40
rect -40 -40 40 40
rect 40 -40 80 40
rect 80 -40 120 40
rect -120 -80 120 -40
rect -120 -120 -80 -80
rect -80 -120 -40 -80
rect -40 -120 40 -80
rect 40 -120 80 -80
rect 80 -120 120 -80
rect 180 -200 420 -180
rect 180 -280 200 -200
rect 200 -280 280 -200
rect 280 -280 420 -200
rect 180 -420 420 -280
<< metal5 >>
tri -861 550 -550 861 se
tri -861 420 -731 550 ne
rect -731 420 -550 550
tri -550 420 -109 861 sw
tri -731 120 -431 420 ne
rect -431 180 -420 420
rect -180 180 -109 420
rect -431 120 -109 180
tri -109 120 191 420 sw
tri -431 -180 -131 120 ne
rect -131 -120 -120 120
rect 120 -120 191 120
rect -131 -180 191 -120
tri 191 -180 491 120 sw
tri -131 -420 109 -180 ne
rect 109 -420 180 -180
rect 420 -420 491 -180
tri 109 -550 239 -420 ne
rect 239 -550 491 -420
tri 491 -550 861 -180 sw
tri 239 -861 550 -550 ne
tri 550 -861 861 -550 nw
<< end >>
