magic
tech sky130A
magscale 1 2
timestamp 1620343632
<< nwell >>
rect -3000 40 3000 4500
<< pwell >>
rect -3000 -4500 3000 -40
<< mvpsubdiff >>
rect -2934 -118 2934 -106
rect -2934 -278 -2700 -118
rect 2700 -278 2934 -118
rect -2934 -290 2934 -278
rect -2934 -340 -2750 -290
rect -2934 -4200 -2922 -340
rect -2762 -4200 -2750 -340
rect -2934 -4250 -2750 -4200
rect 2750 -340 2934 -290
rect 2750 -4200 2762 -340
rect 2922 -4200 2934 -340
rect 2750 -4250 2934 -4200
rect -2934 -4262 2934 -4250
rect -2934 -4422 -2700 -4262
rect 2700 -4422 2934 -4262
rect -2934 -4434 2934 -4422
<< mvnsubdiff >>
rect -2934 4422 2934 4434
rect -2934 4262 -2700 4422
rect 2700 4262 2934 4422
rect -2934 4250 2934 4262
rect -2934 4200 -2750 4250
rect -2934 340 -2922 4200
rect -2762 340 -2750 4200
rect -2934 290 -2750 340
rect 2750 4200 2934 4250
rect 2750 340 2762 4200
rect 2922 340 2934 4200
rect 2750 290 2934 340
rect -2934 278 2934 290
rect -2934 118 -2700 278
rect 2700 118 2934 278
rect -2934 106 2934 118
<< mvpsubdiffcont >>
rect -2700 -278 2700 -118
rect -2922 -4200 -2762 -340
rect 2762 -4200 2922 -340
rect -2700 -4422 2700 -4262
<< mvnsubdiffcont >>
rect -2700 4262 2700 4422
rect -2922 340 -2762 4200
rect 2762 340 2922 4200
rect -2700 118 2700 278
<< locali >>
rect -2922 4200 -2762 4422
rect 2762 4200 2922 4422
rect -1307 2453 -1273 2496
rect -1307 2419 -1227 2453
rect -1227 2245 -1095 2419
rect -969 2345 -837 2419
rect -711 2345 -579 2419
rect -533 2345 -499 2496
rect -453 2345 -321 2419
rect 321 2345 453 2419
rect 499 2345 533 2496
rect 1273 2453 1307 2496
rect 1227 2419 1307 2453
rect 579 2345 711 2419
rect 837 2345 969 2419
rect -969 2285 969 2345
rect 1095 2245 1227 2419
rect -1228 1881 -1095 2245
rect 1094 1881 1227 2245
rect -1228 1821 1227 1881
rect -969 1747 -837 1821
rect -711 1747 -579 1821
rect -453 1747 -321 1821
rect -195 1747 -63 1821
rect 63 1747 195 1821
rect 321 1747 453 1821
rect 579 1747 711 1821
rect 837 1747 969 1821
rect -2922 118 -2762 340
rect 2762 118 2922 340
rect -2922 -340 -2762 -118
rect 2762 -340 2922 -118
rect -969 -588 968 -528
rect -969 -662 -837 -588
rect -711 -662 -579 -588
rect -533 -696 -499 -588
rect -453 -662 -321 -588
rect 321 -662 453 -588
rect 499 -696 533 -588
rect 579 -662 711 -588
rect 837 -662 969 -588
rect -533 -2308 533 -2248
rect -533 -2496 -499 -2308
rect -275 -2388 275 -2348
rect -275 -2496 -241 -2388
rect 241 -2496 275 -2388
rect 499 -2496 533 -2308
rect -2081 -3538 -2047 -3504
rect 2047 -3538 2081 -3504
rect -2081 -3646 -1869 -3538
rect -1485 -3646 -1353 -3538
rect 2001 -3572 2081 -3538
rect -969 -3646 -837 -3572
rect -711 -3646 -579 -3572
rect -453 -3646 -321 -3572
rect -195 -3646 -63 -3572
rect 63 -3646 195 -3572
rect 321 -3646 453 -3572
rect 579 -3646 711 -3572
rect 837 -3646 969 -3572
rect 1353 -3646 1485 -3572
rect 1869 -3646 2081 -3572
rect -2081 -3706 2081 -3646
rect -2922 -4422 -2762 -4200
rect 2762 -4422 2922 -4200
<< viali >>
rect -2762 4262 -2700 4422
rect -2700 4262 2700 4422
rect 2700 4262 2762 4422
rect -2922 477 -2762 4063
rect 2762 477 2922 4063
rect -2762 118 -2700 278
rect -2700 118 2700 278
rect 2700 118 2762 278
rect -2762 -278 -2700 -118
rect -2700 -278 2700 -118
rect 2700 -278 2762 -118
rect -2922 -4063 -2762 -477
rect 2762 -4063 2922 -477
rect -2762 -4422 -2700 -4262
rect -2700 -4422 2700 -4262
rect 2700 -4422 2762 -4262
<< metal1 >>
rect -2928 4422 2928 4428
rect -2928 4262 -2762 4422
rect 2762 4262 2928 4422
rect -2928 4256 2928 4262
rect -2928 4063 -2756 4256
rect -2928 477 -2922 4063
rect -2762 3747 -2756 4063
rect -2156 3956 -2146 4256
rect 2146 3956 2156 4256
rect 2756 4063 2928 4256
rect -539 3837 540 3867
rect -539 3777 -30 3837
rect 30 3777 540 3837
rect -539 3767 540 3777
rect -2762 3627 -1009 3747
rect -2762 1947 -2756 3627
rect -1571 3500 -1525 3627
rect -1465 3541 -1373 3627
rect -1055 3500 -1009 3627
rect -539 3500 -493 3767
rect -175 3685 175 3727
rect -175 3625 -30 3685
rect 30 3625 175 3685
rect -175 3541 175 3625
rect -23 3500 23 3541
rect 493 3500 539 3767
rect 2756 3747 2762 4063
rect 1009 3627 2762 3747
rect 1009 3500 1055 3627
rect 1373 3541 1465 3627
rect 1525 3500 1571 3627
rect -1313 2273 -1267 2500
rect -1217 2346 -1207 2413
rect -1115 2346 -1105 2413
rect -797 2373 -751 2500
rect -281 2373 -235 2500
rect 235 2373 281 2500
rect 751 2373 797 2500
rect -797 2313 797 2373
rect 1267 2273 1313 2500
rect -1313 2213 1313 2273
rect -50 2173 50 2213
rect -1835 2073 -1825 2173
rect -1745 2073 50 2173
rect -2762 1827 -751 1947
rect -2762 477 -2756 1827
rect -1313 1700 -1267 1827
rect -1207 1741 -1115 1827
rect -797 1700 -751 1827
rect -539 1913 539 1959
rect 2756 1947 2762 3627
rect -539 1700 -493 1913
rect -281 1827 281 1873
rect -281 1700 -235 1827
rect 235 1700 281 1827
rect 493 1700 539 1913
rect 751 1827 2762 1947
rect 751 1700 797 1827
rect 1115 1741 1207 1827
rect 1267 1700 1313 1827
rect -1055 573 -1009 700
rect -23 671 23 700
rect -39 613 -29 671
rect 29 613 39 671
rect 1009 573 1055 700
rect -1055 513 1055 573
rect -2928 284 -2756 477
rect -30 468 30 513
rect 2756 477 2762 1827
rect 2922 477 2928 4063
rect -40 408 -30 468
rect 30 408 40 468
rect 2756 284 2928 477
rect -2928 278 2928 284
rect -2928 118 -2762 278
rect 2762 118 2928 278
rect -2928 112 2928 118
rect -2928 -118 2928 -112
rect -2928 -278 -2762 -118
rect 2762 -278 2928 -118
rect -2928 -284 2928 -278
rect -2928 -477 -2756 -284
rect -2928 -4063 -2922 -477
rect -2762 -1827 -2756 -477
rect -39 -409 75 -349
rect 135 -409 145 -349
rect -39 -513 39 -409
rect 2756 -477 2928 -284
rect -539 -573 539 -513
rect -539 -700 -493 -573
rect -175 -680 -29 -622
rect 29 -680 175 -622
rect -23 -700 23 -680
rect 493 -700 539 -573
rect -1313 -1827 -1267 -1700
rect -1207 -1827 -1115 -1732
rect -1055 -1827 -1009 -1700
rect -2762 -1927 -1009 -1827
rect -797 -1827 -751 -1700
rect -281 -1827 -235 -1700
rect 235 -1827 281 -1700
rect 751 -1827 797 -1700
rect -797 -1927 797 -1827
rect 1009 -1827 1055 -1700
rect 1115 -1827 1207 -1732
rect 1267 -1827 1313 -1700
rect 2756 -1827 2762 -477
rect 1009 -1927 2762 -1827
rect -2762 -2273 -2756 -1927
rect -40 -2210 -30 -2150
rect 30 -2210 40 -2150
rect -2762 -2373 -751 -2273
rect -2762 -4063 -2756 -2373
rect -2345 -2500 -2299 -2373
rect -2239 -2468 -2147 -2373
rect -1829 -2500 -1783 -2373
rect -1723 -2468 -1631 -2373
rect -1313 -2500 -1267 -2373
rect -1207 -2468 -1115 -2373
rect -1072 -2480 -1062 -2420
rect -1002 -2480 -992 -2420
rect -1055 -2500 -1009 -2480
rect -797 -2500 -751 -2373
rect -23 -2500 23 -2210
rect 2756 -2273 2762 -1927
rect 751 -2373 2762 -2273
rect 751 -2500 797 -2373
rect 992 -2480 1002 -2420
rect 1062 -2480 1072 -2420
rect 1115 -2468 1207 -2373
rect 1009 -2500 1055 -2480
rect 1267 -2500 1313 -2373
rect 1631 -2468 1723 -2373
rect 1783 -2500 1829 -2373
rect 2147 -2468 2239 -2373
rect 2299 -2500 2345 -2373
rect -2087 -3728 -2041 -3500
rect -1981 -3546 -1889 -3532
rect -1991 -3606 -1981 -3546
rect -1889 -3606 -1879 -3546
rect -1981 -3728 -1889 -3606
rect -1571 -3668 -1525 -3500
rect 1525 -3668 1571 -3500
rect -1571 -3701 1571 -3668
rect -2087 -3828 -1632 -3728
rect -1571 -3761 -30 -3701
rect 30 -3761 1571 -3701
rect 1889 -3728 1981 -3532
rect 2041 -3728 2087 -3500
rect -1571 -3788 1571 -3761
rect 1632 -3828 2087 -3728
rect -2087 -3846 2087 -3828
rect -2087 -3926 -39 -3846
rect 41 -3926 2087 -3846
rect -2087 -3948 2087 -3926
rect -2928 -4256 -2756 -4063
rect -2156 -4256 -2146 -3956
rect 2146 -4256 2156 -3956
rect 2756 -4063 2762 -2373
rect 2922 -4063 2928 -477
rect 2756 -4256 2928 -4063
rect -2928 -4262 2928 -4256
rect -2928 -4422 -2762 -4262
rect 2762 -4422 2928 -4262
rect -2928 -4428 2928 -4422
<< via1 >>
rect -2756 3956 -2156 4256
rect 2156 3956 2756 4256
rect -30 3777 30 3837
rect -30 3625 30 3685
rect -1207 2346 -1115 2413
rect -1825 2073 -1745 2173
rect -29 613 29 671
rect -30 408 30 468
rect 75 -409 135 -349
rect -29 -680 29 -622
rect -30 -2210 30 -2150
rect -1062 -2480 -1002 -2420
rect 1002 -2480 1062 -2420
rect -1981 -3606 -1889 -3546
rect -30 -3761 30 -3701
rect -39 -3926 41 -3846
rect -2756 -4256 -2156 -3956
rect 2156 -4256 2756 -3956
<< metal2 >>
rect -2756 4256 -2156 4266
rect -2756 3946 -2156 3956
rect 2156 4256 2756 4266
rect 2156 3946 2756 3956
rect -30 3837 1884 3887
rect 30 3777 1884 3837
rect -30 3767 1884 3777
rect -1683 3685 1695 3695
rect -1683 3625 -30 3685
rect 30 3625 1695 3685
rect -1683 3616 1695 3625
rect -1683 3615 30 3616
rect -1683 2187 -1603 3615
rect -1207 2413 -1115 2423
rect -1207 2336 -1115 2346
rect -1865 2173 -1745 2183
rect -1865 2073 -1825 2173
rect -1683 2097 -1603 2107
rect -1865 -2184 -1745 2073
rect -29 671 29 681
rect -29 597 29 613
rect -29 519 170 597
rect -70 468 30 478
rect -70 408 -30 468
rect -70 -498 30 408
rect 70 -349 170 519
rect 70 -409 75 -349
rect 135 -409 170 -349
rect 70 -419 170 -409
rect -70 -508 40 -498
rect -70 -588 -40 -508
rect -70 -598 40 -588
rect -30 -622 30 -598
rect -30 -680 -29 -622
rect 29 -680 30 -622
rect -30 -690 30 -680
rect 1575 -1982 1695 3616
rect -2537 -2264 -1745 -2184
rect -176 -2061 1695 -1982
rect -176 -2241 -97 -2061
rect 1764 -2140 1884 3767
rect -30 -2150 1884 -2140
rect 30 -2210 1884 -2150
rect -30 -2220 1884 -2210
rect -2537 -3691 -2457 -2264
rect -177 -2350 -96 -2241
rect -30 -2350 30 -2348
rect -1062 -2410 1062 -2350
rect -1062 -2420 -1002 -2410
rect -1062 -2490 -1002 -2480
rect 1002 -2420 1062 -2410
rect 1002 -2490 1062 -2480
rect -2269 -3536 -2189 -3526
rect -2189 -3616 -2073 -3536
rect -1981 -3546 -1889 -3536
rect -1981 -3616 -1889 -3606
rect -2269 -3626 -2189 -3616
rect -2537 -3701 30 -3691
rect -2537 -3761 -30 -3701
rect -2537 -3771 30 -3761
rect -39 -3846 41 -3836
rect -39 -3936 41 -3926
rect -2756 -3956 -2156 -3946
rect -2756 -4266 -2156 -4256
rect 2156 -3956 2756 -3946
rect 2156 -4266 2756 -4256
<< rmetal2 >>
rect -2073 -3616 -1981 -3536
<< via2 >>
rect -2756 3956 -2156 4256
rect 2156 3956 2756 4256
rect -1207 2346 -1115 2413
rect -1683 2107 -1603 2187
rect -40 -588 40 -508
rect -2269 -3616 -2189 -3536
rect -39 -3926 41 -3846
rect -2756 -4256 -2156 -3956
rect 2156 -4256 2756 -3956
<< metal3 >>
rect -2766 4256 -2146 4261
rect -2766 3956 -2756 4256
rect -2156 3956 -2146 4256
rect -2766 3951 -2146 3956
rect 2146 4256 2766 4261
rect 2146 3956 2156 4256
rect 2756 3956 2766 4256
rect 2146 3951 2766 3956
rect -2641 2413 -1105 2418
rect -2641 2346 -1207 2413
rect -1115 2346 -1105 2413
rect -2641 2318 -1105 2346
rect -1693 2187 -1593 2192
rect -2641 2107 -1683 2187
rect -1603 2107 -1593 2187
rect -2641 2087 -1593 2107
rect -2641 -508 50 -480
rect -2641 -580 -40 -508
rect -50 -588 -40 -580
rect 40 -588 50 -508
rect -50 -593 50 -588
rect -2641 -824 -2325 -734
rect -2641 -2862 -2500 -2742
rect -2589 -3124 -2500 -2862
rect -2590 -3710 -2500 -3124
rect -2415 -3531 -2325 -824
rect -2415 -3536 -2179 -3531
rect -2415 -3616 -2269 -3536
rect -2189 -3616 -2179 -3536
rect -2415 -3621 -2179 -3616
rect -2590 -3800 -1674 -3710
rect -1764 -3841 -1674 -3800
rect -1764 -3846 51 -3841
rect -1764 -3926 -39 -3846
rect 41 -3926 51 -3846
rect -1764 -3931 51 -3926
rect -2766 -3956 -2146 -3951
rect -2766 -4256 -2756 -3956
rect -2156 -4256 -2146 -3956
rect -2766 -4261 -2146 -4256
rect 2146 -3956 2766 -3951
rect 2146 -4256 2156 -3956
rect 2756 -4256 2766 -3956
rect 2146 -4261 2766 -4256
<< via3 >>
rect -2756 3956 -2156 4256
rect 2156 3956 2756 4256
rect -2756 -4256 -2156 -3956
rect 2156 -4256 2756 -3956
<< metal4 >>
rect -3000 4256 3000 4500
rect -3000 3956 -2756 4256
rect -2156 3956 2156 4256
rect 2756 3956 3000 4256
rect -3000 3700 3000 3956
rect -3000 -3956 3000 -3700
rect -3000 -4256 -2756 -3956
rect -2156 -4256 2156 -3956
rect 2756 -4256 3000 -3956
rect -3000 -4500 3000 -4256
use sky130_fd_pr__nfet_g5v0d10v5_V2YKKA  xm1
timestamp 1620252470
transform 1 0 0 0 1 -1200
box -1319 -588 1319 588
use sky130_fd_pr__nfet_g5v0d10v5_7QEKRB  xm2
timestamp 1620252470
transform 1 0 0 0 1 -3000
box -2351 -588 2351 588
use sky130_fd_pr__pfet_g5v0d10v5_QRGZLW  xm3
timestamp 1620252470
transform 1 0 0 0 1 1200
box -1385 -600 1385 600
use sky130_fd_pr__pfet_g5v0d10v5_QNH2MW  xm4
timestamp 1620252470
transform 1 0 0 0 1 3000
box -1643 -600 1643 600
<< labels >>
flabel metal4 -3000 3700 -3000 4500 3 FreeSans 480 0 0 0 vdd
port 1 e
flabel metal4 -3000 -4500 -3000 -3700 3 FreeSans 480 0 0 0 vss
port 2 e
flabel metal3 -2641 -580 -2641 -480 1 FreeSans 240 0 0 0 vcn
port 3 n
flabel metal3 -2641 2087 -2641 2187 1 FreeSans 240 0 0 0 vcp
port 4 n
flabel metal3 -2641 2318 -2641 2418 1 FreeSans 240 0 0 0 vbp
port 5 n
flabel metal3 -2641 -824 -2641 -734 1 FreeSans 240 0 0 0 vbn
port 6 n
flabel metal3 -2641 -2862 -2641 -2742 1 FreeSans 240 0 0 0 ibias
port 7 n
<< properties >>
string FIXED_BBOX -2842 -4342 2842 -198
<< end >>
